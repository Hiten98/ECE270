// 4 bit ring counter
module ring_counter(CLK, R, Q);
  begin
  end
