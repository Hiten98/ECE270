module button( );


endmodule

