module selfCorrecting_johnson_counter(CLK, R, Q);
