// 4 bit ring counter
module ring_counter(CLK, R, Q);
  begin
  always @ (posedge CLK)
    begin
    end
  end
